`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2019/04/12 12:25:00
// Design Name: 
// Module Name: signal_process
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module signal_process(
    input [3:0]dir_shake_removed,
    input clk_100M,
    output 
);
   
   
   
   
   
   
   
   
   
   
   
   /* localparam S0=2'b00,S1=2'b01,S2=2'b10;
    reg [1:0]state=S0;
    
	always@(posedge clk_100M) 
	begin
	   case(state)
	   S0: if(in)  state<=S1;
	       else    state<=S0;
	   S1: if(in)  state<=S2;
	       else    state<=S0;
	   S2: if(in)  state<=S2;
	       else    state<=S0;
	   endcase
    end
    
    always @(state)
    begin
        case(state)
        S0: out = 0;
        S1: out = 1;
        S2: out = 0;
        endcase
    end*/
endmodule
